module Mux12bit_12(p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,address,Dout);

input [11:0] p0;
input [11:0] p1;
input [11:0] p2;
input [11:0] p3;
input [11:0] p4;
input [11:0] p5;
input [11:0] p6;
input [11:0] p7;
input [11:0] p8;
input [11:0] p9;
input [11:0] p10;
input [11:0] p11;
input [3:0] address;
output [11:0] Dout;

wire [11:0] b131;
wire [11:0] b122;
wire [11:0] b130;
wire [11:0] b129;
wire [11:0] b128;
wire [11:0] b127;
wire [11:0] b126;
wire [11:0] b125;
wire [11:0] b124;
wire [11:0] b123;
wire [11:0] b121;
wire [11:0] b120;
wire [3:0] b156;
wire [11:0] b164;
wire  b131_0_w12;
wire  b122_0_w13;
wire  b130_0_w14;
wire  b129_0_w15;
wire  b128_0_w16;
wire  b127_0_w17;
wire  b126_0_w18;
wire  b125_0_w19;
wire  b124_0_w20;
wire  b123_0_w21;
wire  b121_0_w22;
wire  b120_0_w23;
wire  b131_1_w25;
wire  b122_1_w26;
wire  b130_1_w27;
wire  b129_1_w28;
wire  b128_1_w29;
wire  b127_1_w30;
wire  b126_1_w31;
wire  b125_1_w32;
wire  b124_1_w33;
wire  b123_1_w34;
wire  b121_1_w35;
wire  b120_1_w36;
wire  b131_2_w37;
wire  b122_2_w38;
wire  b130_2_w39;
wire  b129_2_w40;
wire  b128_2_w41;
wire  b127_2_w42;
wire  b126_2_w43;
wire  b125_2_w44;
wire  b124_2_w45;
wire  b123_2_w46;
wire  b121_2_w47;
wire  b120_2_w48;
wire  b131_3_w49;
wire  b122_3_w50;
wire  b130_3_w51;
wire  b129_3_w52;
wire  b128_3_w53;
wire  b127_3_w54;
wire  b126_3_w55;
wire  b125_3_w56;
wire  b124_3_w57;
wire  b123_3_w58;
wire  b121_3_w59;
wire  b120_3_w60;
wire  b131_4_w61;
wire  b122_4_w62;
wire  b130_4_w63;
wire  b129_4_w64;
wire  b128_4_w65;
wire  b127_4_w66;
wire  b126_4_w67;
wire  b125_4_w68;
wire  b124_4_w69;
wire  b123_4_w70;
wire  b121_4_w71;
wire  b120_4_w72;
wire  b131_5_w73;
wire  b122_5_w74;
wire  b130_5_w75;
wire  b129_5_w76;
wire  b128_5_w77;
wire  b127_5_w78;
wire  b126_5_w79;
wire  b125_5_w80;
wire  b124_5_w81;
wire  b123_5_w82;
wire  b121_5_w83;
wire  b120_5_w84;
wire  b131_6_w85;
wire  b122_6_w86;
wire  b130_6_w87;
wire  b129_6_w88;
wire  b128_6_w89;
wire  b127_6_w90;
wire  b126_6_w91;
wire  b125_6_w92;
wire  b124_6_w93;
wire  b123_6_w94;
wire  b121_6_w95;
wire  b120_6_w96;
wire  b131_7_w97;
wire  b122_7_w98;
wire  b130_7_w99;
wire  b129_7_w100;
wire  b128_7_w101;
wire  b127_7_w102;
wire  b126_7_w103;
wire  b125_7_w104;
wire  b124_7_w105;
wire  b123_7_w106;
wire  b121_7_w107;
wire  b120_7_w108;
wire  b131_8_w109;
wire  b122_8_w110;
wire  b130_8_w111;
wire  b129_8_w112;
wire  b128_8_w113;
wire  b127_8_w114;
wire  b126_8_w115;
wire  b125_8_w116;
wire  b124_8_w117;
wire  b123_8_w118;
wire  b121_8_w119;
wire  b120_8_w120;
wire  b131_9_w121;
wire  b122_9_w122;
wire  b130_9_w123;
wire  b129_9_w124;
wire  b128_9_w125;
wire  b127_9_w126;
wire  b126_9_w127;
wire  b125_9_w128;
wire  b124_9_w129;
wire  b123_9_w130;
wire  b121_9_w131;
wire  b120_9_w132;
wire  b131_10_w133;
wire  b122_10_w134;
wire  b130_10_w135;
wire  b129_10_w136;
wire  b128_10_w137;
wire  b127_10_w138;
wire  b126_10_w139;
wire  b125_10_w140;
wire  b124_10_w141;
wire  b123_10_w142;
wire  b121_10_w143;
wire  b120_10_w144;
wire  b131_11_w145;
wire  b122_11_w146;
wire  b130_11_w147;
wire  b129_11_w148;
wire  b128_11_w149;
wire  b127_11_w150;
wire  b126_11_w151;
wire  b125_11_w152;
wire  b124_11_w153;
wire  b123_11_w154;
wire  b121_11_w155;
wire  b120_11_w156;
wire  b164_0;
wire  b164_1;
wire  b164_2;
wire  b164_3;
wire  b164_4;
wire  b164_5;
wire  b164_6;
wire  b164_7;
wire  b164_8;
wire  b164_9;
wire  b164_10;
wire  b164_11;

assign b131 = p0;
assign b130 = p1;
assign b129 = p2;
assign b128 = p3;
assign b127 = p4;
assign b126 = p5;
assign b125 = p6;
assign b124 = p7;
assign b123 = p8;
assign b122 = p9;
assign b121 = p10;
assign b120 = p11;
assign b156 = address;
assign Dout = b164;

assign b164[11] = b164_11;
assign b164[10] = b164_10;
assign b164[9] = b164_9;
assign b164[8] = b164_8;
assign b164[7] = b164_7;
assign b164[6] = b164_6;
assign b164[5] = b164_5;
assign b164[4] = b164_4;
assign b164[3] = b164_3;
assign b164[2] = b164_2;
assign b164[1] = b164_1;
assign b164[0] = b164_0;

assign b131_0_w12 = {b131[0]};
assign b122_0_w13 = {b122[0]};
assign b130_0_w14 = {b130[0]};
assign b129_0_w15 = {b129[0]};
assign b128_0_w16 = {b128[0]};
assign b127_0_w17 = {b127[0]};
assign b126_0_w18 = {b126[0]};
assign b125_0_w19 = {b125[0]};
assign b124_0_w20 = {b124[0]};
assign b123_0_w21 = {b123[0]};
assign b121_0_w22 = {b121[0]};
assign b120_0_w23 = {b120[0]};
assign b131_1_w25 = {b131[1]};
assign b122_1_w26 = {b122[1]};
assign b130_1_w27 = {b130[1]};
assign b129_1_w28 = {b129[1]};
assign b128_1_w29 = {b128[1]};
assign b127_1_w30 = {b127[1]};
assign b126_1_w31 = {b126[1]};
assign b125_1_w32 = {b125[1]};
assign b124_1_w33 = {b124[1]};
assign b123_1_w34 = {b123[1]};
assign b121_1_w35 = {b121[1]};
assign b120_1_w36 = {b120[1]};
assign b131_2_w37 = {b131[2]};
assign b122_2_w38 = {b122[2]};
assign b130_2_w39 = {b130[2]};
assign b129_2_w40 = {b129[2]};
assign b128_2_w41 = {b128[2]};
assign b127_2_w42 = {b127[2]};
assign b126_2_w43 = {b126[2]};
assign b125_2_w44 = {b125[2]};
assign b124_2_w45 = {b124[2]};
assign b123_2_w46 = {b123[2]};
assign b121_2_w47 = {b121[2]};
assign b120_2_w48 = {b120[2]};
assign b131_3_w49 = {b131[3]};
assign b122_3_w50 = {b122[3]};
assign b130_3_w51 = {b130[3]};
assign b129_3_w52 = {b129[3]};
assign b128_3_w53 = {b128[3]};
assign b127_3_w54 = {b127[3]};
assign b126_3_w55 = {b126[3]};
assign b125_3_w56 = {b125[3]};
assign b124_3_w57 = {b124[3]};
assign b123_3_w58 = {b123[3]};
assign b121_3_w59 = {b121[3]};
assign b120_3_w60 = {b120[3]};
assign b131_4_w61 = {b131[4]};
assign b122_4_w62 = {b122[4]};
assign b130_4_w63 = {b130[4]};
assign b129_4_w64 = {b129[4]};
assign b128_4_w65 = {b128[4]};
assign b127_4_w66 = {b127[4]};
assign b126_4_w67 = {b126[4]};
assign b125_4_w68 = {b125[4]};
assign b124_4_w69 = {b124[4]};
assign b123_4_w70 = {b123[4]};
assign b121_4_w71 = {b121[4]};
assign b120_4_w72 = {b120[4]};
assign b131_5_w73 = {b131[5]};
assign b122_5_w74 = {b122[5]};
assign b130_5_w75 = {b130[5]};
assign b129_5_w76 = {b129[5]};
assign b128_5_w77 = {b128[5]};
assign b127_5_w78 = {b127[5]};
assign b126_5_w79 = {b126[5]};
assign b125_5_w80 = {b125[5]};
assign b124_5_w81 = {b124[5]};
assign b123_5_w82 = {b123[5]};
assign b121_5_w83 = {b121[5]};
assign b120_5_w84 = {b120[5]};
assign b131_6_w85 = {b131[6]};
assign b122_6_w86 = {b122[6]};
assign b130_6_w87 = {b130[6]};
assign b129_6_w88 = {b129[6]};
assign b128_6_w89 = {b128[6]};
assign b127_6_w90 = {b127[6]};
assign b126_6_w91 = {b126[6]};
assign b125_6_w92 = {b125[6]};
assign b124_6_w93 = {b124[6]};
assign b123_6_w94 = {b123[6]};
assign b121_6_w95 = {b121[6]};
assign b120_6_w96 = {b120[6]};
assign b131_7_w97 = {b131[7]};
assign b122_7_w98 = {b122[7]};
assign b130_7_w99 = {b130[7]};
assign b129_7_w100 = {b129[7]};
assign b128_7_w101 = {b128[7]};
assign b127_7_w102 = {b127[7]};
assign b126_7_w103 = {b126[7]};
assign b125_7_w104 = {b125[7]};
assign b124_7_w105 = {b124[7]};
assign b123_7_w106 = {b123[7]};
assign b121_7_w107 = {b121[7]};
assign b120_7_w108 = {b120[7]};
assign b131_8_w109 = {b131[8]};
assign b122_8_w110 = {b122[8]};
assign b130_8_w111 = {b130[8]};
assign b129_8_w112 = {b129[8]};
assign b128_8_w113 = {b128[8]};
assign b127_8_w114 = {b127[8]};
assign b126_8_w115 = {b126[8]};
assign b125_8_w116 = {b125[8]};
assign b124_8_w117 = {b124[8]};
assign b123_8_w118 = {b123[8]};
assign b121_8_w119 = {b121[8]};
assign b120_8_w120 = {b120[8]};
assign b131_9_w121 = {b131[9]};
assign b122_9_w122 = {b122[9]};
assign b130_9_w123 = {b130[9]};
assign b129_9_w124 = {b129[9]};
assign b128_9_w125 = {b128[9]};
assign b127_9_w126 = {b127[9]};
assign b126_9_w127 = {b126[9]};
assign b125_9_w128 = {b125[9]};
assign b124_9_w129 = {b124[9]};
assign b123_9_w130 = {b123[9]};
assign b121_9_w131 = {b121[9]};
assign b120_9_w132 = {b120[9]};
assign b131_10_w133 = {b131[10]};
assign b122_10_w134 = {b122[10]};
assign b130_10_w135 = {b130[10]};
assign b129_10_w136 = {b129[10]};
assign b128_10_w137 = {b128[10]};
assign b127_10_w138 = {b127[10]};
assign b126_10_w139 = {b126[10]};
assign b125_10_w140 = {b125[10]};
assign b124_10_w141 = {b124[10]};
assign b123_10_w142 = {b123[10]};
assign b121_10_w143 = {b121[10]};
assign b120_10_w144 = {b120[10]};
assign b131_11_w145 = {b131[11]};
assign b122_11_w146 = {b122[11]};
assign b130_11_w147 = {b130[11]};
assign b129_11_w148 = {b129[11]};
assign b128_11_w149 = {b128[11]};
assign b127_11_w150 = {b127[11]};
assign b126_11_w151 = {b126[11]};
assign b125_11_w152 = {b125[11]};
assign b124_11_w153 = {b124[11]};
assign b123_11_w154 = {b123[11]};
assign b121_11_w155 = {b121[11]};
assign b120_11_w156 = {b120[11]};

Mux12bit_4
     s0 (
      .D1(b131_0_w12),
      .D0(b122_0_w13),
      .D2(b130_0_w14),
      .D3(b129_0_w15),
      .D4(b128_0_w16),
      .D5(b127_0_w17),
      .D6(b126_0_w18),
      .D7(b125_0_w19),
      .D8(b124_0_w20),
      .D9(b123_0_w21),
      .D_sharp(b121_0_w22),
      .D_star(b120_0_w23),
      .B_in(b156),
      .D_out(b164_0));

Mux12bit_4
     s1 (
      .D1(b131_1_w25),
      .D0(b122_1_w26),
      .D2(b130_1_w27),
      .D3(b129_1_w28),
      .D4(b128_1_w29),
      .D5(b127_1_w30),
      .D6(b126_1_w31),
      .D7(b125_1_w32),
      .D8(b124_1_w33),
      .D9(b123_1_w34),
      .D_sharp(b121_1_w35),
      .D_star(b120_1_w36),
      .B_in(b156),
      .D_out(b164_1));

Mux12bit_4
     s2 (
      .D1(b131_2_w37),
      .D0(b122_2_w38),
      .D2(b130_2_w39),
      .D3(b129_2_w40),
      .D4(b128_2_w41),
      .D5(b127_2_w42),
      .D6(b126_2_w43),
      .D7(b125_2_w44),
      .D8(b124_2_w45),
      .D9(b123_2_w46),
      .D_sharp(b121_2_w47),
      .D_star(b120_2_w48),
      .B_in(b156),
      .D_out(b164_2));

Mux12bit_4
     s3 (
      .D1(b131_3_w49),
      .D0(b122_3_w50),
      .D2(b130_3_w51),
      .D3(b129_3_w52),
      .D4(b128_3_w53),
      .D5(b127_3_w54),
      .D6(b126_3_w55),
      .D7(b125_3_w56),
      .D8(b124_3_w57),
      .D9(b123_3_w58),
      .D_sharp(b121_3_w59),
      .D_star(b120_3_w60),
      .B_in(b156),
      .D_out(b164_3));

Mux12bit_4
     s4 (
      .D1(b131_4_w61),
      .D0(b122_4_w62),
      .D2(b130_4_w63),
      .D3(b129_4_w64),
      .D4(b128_4_w65),
      .D5(b127_4_w66),
      .D6(b126_4_w67),
      .D7(b125_4_w68),
      .D8(b124_4_w69),
      .D9(b123_4_w70),
      .D_sharp(b121_4_w71),
      .D_star(b120_4_w72),
      .B_in(b156),
      .D_out(b164_4));

Mux12bit_4
     s5 (
      .D1(b131_5_w73),
      .D0(b122_5_w74),
      .D2(b130_5_w75),
      .D3(b129_5_w76),
      .D4(b128_5_w77),
      .D5(b127_5_w78),
      .D6(b126_5_w79),
      .D7(b125_5_w80),
      .D8(b124_5_w81),
      .D9(b123_5_w82),
      .D_sharp(b121_5_w83),
      .D_star(b120_5_w84),
      .B_in(b156),
      .D_out(b164_5));

Mux12bit_4
     s6 (
      .D1(b131_6_w85),
      .D0(b122_6_w86),
      .D2(b130_6_w87),
      .D3(b129_6_w88),
      .D4(b128_6_w89),
      .D5(b127_6_w90),
      .D6(b126_6_w91),
      .D7(b125_6_w92),
      .D8(b124_6_w93),
      .D9(b123_6_w94),
      .D_sharp(b121_6_w95),
      .D_star(b120_6_w96),
      .B_in(b156),
      .D_out(b164_6));

Mux12bit_4
     s7 (
      .D1(b131_7_w97),
      .D0(b122_7_w98),
      .D2(b130_7_w99),
      .D3(b129_7_w100),
      .D4(b128_7_w101),
      .D5(b127_7_w102),
      .D6(b126_7_w103),
      .D7(b125_7_w104),
      .D8(b124_7_w105),
      .D9(b123_7_w106),
      .D_sharp(b121_7_w107),
      .D_star(b120_7_w108),
      .B_in(b156),
      .D_out(b164_7));

Mux12bit_4
     s8 (
      .D1(b131_8_w109),
      .D0(b122_8_w110),
      .D2(b130_8_w111),
      .D3(b129_8_w112),
      .D4(b128_8_w113),
      .D5(b127_8_w114),
      .D6(b126_8_w115),
      .D7(b125_8_w116),
      .D8(b124_8_w117),
      .D9(b123_8_w118),
      .D_sharp(b121_8_w119),
      .D_star(b120_8_w120),
      .B_in(b156),
      .D_out(b164_8));

Mux12bit_4
     s9 (
      .D1(b131_9_w121),
      .D0(b122_9_w122),
      .D2(b130_9_w123),
      .D3(b129_9_w124),
      .D4(b128_9_w125),
      .D5(b127_9_w126),
      .D6(b126_9_w127),
      .D7(b125_9_w128),
      .D8(b124_9_w129),
      .D9(b123_9_w130),
      .D_sharp(b121_9_w131),
      .D_star(b120_9_w132),
      .B_in(b156),
      .D_out(b164_9));

Mux12bit_4
     s10 (
      .D1(b131_10_w133),
      .D0(b122_10_w134),
      .D2(b130_10_w135),
      .D3(b129_10_w136),
      .D4(b128_10_w137),
      .D5(b127_10_w138),
      .D6(b126_10_w139),
      .D7(b125_10_w140),
      .D8(b124_10_w141),
      .D9(b123_10_w142),
      .D_sharp(b121_10_w143),
      .D_star(b120_10_w144),
      .B_in(b156),
      .D_out(b164_10));

Mux12bit_4
     s11 (
      .D1(b131_11_w145),
      .D0(b122_11_w146),
      .D2(b130_11_w147),
      .D3(b129_11_w148),
      .D4(b128_11_w149),
      .D5(b127_11_w150),
      .D6(b126_11_w151),
      .D7(b125_11_w152),
      .D8(b124_11_w153),
      .D9(b123_11_w154),
      .D_sharp(b121_11_w155),
      .D_star(b120_11_w156),
      .B_in(b156),
      .D_out(b164_11));

endmodule

