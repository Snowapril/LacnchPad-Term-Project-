module MUX4bit_4_tb;

reg [3:0] D0;
reg [3:0] D1;
reg [3:0] D2;
reg [3:0] D3;
wire [3:0] Dout;
reg S0;
reg S1;

MUX4bit_4
 U0 (
  .D0(D0),
  .D1(D1),
  .D2(D2),
  .D3(D3),
  .Dout(Dout),
  .S0(S0),
  .S1(S1));

  initial
  begin
    D0 = 4'b1010;
    #200 D0 = 4'b1111;
    #400 D0 = 4'b1001;
    #200 D0 = 4'b0110;
    #200 D0 = 4'b1110;
    #200 D0 = 4'b0010;
    #200 D0 = 4'b1111;
    #200 D0 = 4'b0001;
    #200 D0 = 4'b1011;
    #200 D0 = 4'b1000;
    #400 D0 = 4'b0000;
    #400 D0 = 4'b1001;
    #200 D0 = 4'b0000;
    #200 D0 = 4'b1001;
    #200 D0 = 4'b1010;
    #200 D0 = 4'b0011;
    #200 D0 = 4'b1010;
    #200 D0 = 4'b0011;
    #200 D0 = 4'b0010;
    #200 D0 = 4'b0111;
    #600 D0 = 4'b0011;
    #200 D0 = 4'b1000;
    #200 D0 = 4'b1001;
    #200 D0 = 4'b1100;
    #200 D0 = 4'b0100;
    #200 D0 = 4'b0010;
    #200 D0 = 4'b1010;
    #200 D0 = 4'b0110;
    #200 D0 = 4'b1011;
    #200 D0 = 4'b0010;
    #200 D0 = 4'b1111;
    #200 D0 = 4'b1011;
    #200 D0 = 4'b0000;
    #200 D0 = 4'b0010;
    #200 D0 = 4'b0100;
    #200 D0 = 4'b0010;
    #400 D0 = 4'b0111;
    #400 D0 = 4'b0001;
    #200 D0 = 4'b0000;
    #200 D0 = 4'b1100;
    #200 D0 = 4'b1011;
    #200 D0 = 4'b1010;
    #200 D0 = 4'b1001;
  end

  initial
  begin
    D1 = 4'b1001;
    #200 D1 = 4'b1000;
    #200 D1 = 4'b0110;
    #200 D1 = 4'b1101;
    #200 D1 = 4'b1011;
    #200 D1 = 4'b1100;
    #200 D1 = 4'b0111;
    #200 D1 = 4'b0010;
    #400 D1 = 4'b1010;
    #200 D1 = 4'b1111;
    #200 D1 = 4'b0000;
    #200 D1 = 4'b1110;
    #200 D1 = 4'b1011;
    #200 D1 = 4'b0010;
    #200 D1 = 4'b1100;
    #200 D1 = 4'b1001;
    #200 D1 = 4'b0110;
    #400 D1 = 4'b0101;
    #200 D1 = 4'b1100;
    #200 D1 = 4'b0100;
    #200 D1 = 4'b0101;
    #200 D1 = 4'b1111;
    #200 D1 = 4'b0110;
    #200 D1 = 4'b0000;
    #200 D1 = 4'b1110;
    #200 D1 = 4'b1100;
    #200 D1 = 4'b1011;
    #200 D1 = 4'b0101;
    #200 D1 = 4'b1001;
    #200 D1 = 4'b0110;
    #200 D1 = 4'b0111;
    #200 D1 = 4'b0011;
    #200 D1 = 4'b1001;
    #600 D1 = 4'b0011;
    #200 D1 = 4'b1001;
    #200 D1 = 4'b0100;
    #200 D1 = 4'b1010;
    #200 D1 = 4'b0000;
    #200 D1 = 4'b1011;
    #200 D1 = 4'b1010;
    #400 D1 = 4'b0110;
    #200 D1 = 4'b0011;
    #200 D1 = 4'b1100;
    #200 D1 = 4'b0101;
    #200 D1 = 4'b1111;
  end

  initial
  begin
    D2 = 4'b1000;
    #200 D2 = 4'b0010;
    #400 D2 = 4'b1111;
    #200 D2 = 4'b1110;
    #200 D2 = 4'b0001;
    #200 D2 = 4'b0011;
    #200 D2 = 4'b1001;
    #200 D2 = 4'b1110;
    #200 D2 = 4'b1100;
    #200 D2 = 4'b1000;
    #200 D2 = 4'b1110;
    #200 D2 = 4'b0111;
    #200 D2 = 4'b0000;
    #200 D2 = 4'b0010;
    #200 D2 = 4'b1000;
    #200 D2 = 4'b0111;
    #200 D2 = 4'b0010;
    #200 D2 = 4'b1101;
    #200 D2 = 4'b1010;
    #200 D2 = 4'b1000;
    #200 D2 = 4'b1100;
    #200 D2 = 4'b1111;
    #200 D2 = 4'b1010;
    #200 D2 = 4'b1110;
    #200 D2 = 4'b1010;
    #200 D2 = 4'b1100;
    #200 D2 = 4'b0111;
    #200 D2 = 4'b0100;
    #200 D2 = 4'b1001;
    #200 D2 = 4'b0010;
    #200 D2 = 4'b0000;
    #200 D2 = 4'b1001;
    #200 D2 = 4'b1000;
    #200 D2 = 4'b0011;
    #200 D2 = 4'b1100;
    #200 D2 = 4'b1001;
    #200 D2 = 4'b1011;
    #200 D2 = 4'b1000;
    #200 D2 = 4'b0001;
    #200 D2 = 4'b1110;
    #200 D2 = 4'b0100;
    #200 D2 = 4'b0010;
    #200 D2 = 4'b0110;
    #200 D2 = 4'b0101;
    #200 D2 = 4'b0100;
    #200 D2 = 4'b0011;
    #200 D2 = 4'b0010;
    #200 D2 = 4'b1001;
    #200 D2 = 4'b0100;
  end

  initial
  begin
    D3 = 4'b1000;
    #200 D3 = 4'b0001;
    #200 D3 = 4'b0111;
    #200 D3 = 4'b1101;
    #400 D3 = 4'b1100;
    #200 D3 = 4'b1010;
    #200 D3 = 4'b1110;
    #200 D3 = 4'b0100;
    #200 D3 = 4'b1101;
    #200 D3 = 4'b1001;
    #200 D3 = 4'b1101;
    #200 D3 = 4'b0111;
    #200 D3 = 4'b0110;
    #200 D3 = 4'b0011;
    #200 D3 = 4'b0001;
    #200 D3 = 4'b0100;
    #200 D3 = 4'b1001;
    #200 D3 = 4'b0100;
    #200 D3 = 4'b0001;
    #200 D3 = 4'b0011;
    #200 D3 = 4'b1011;
    #200 D3 = 4'b1100;
    #200 D3 = 4'b0011;
    #200 D3 = 4'b1001;
    #200 D3 = 4'b0000;
    #200 D3 = 4'b1011;
    #200 D3 = 4'b0101;
    #200 D3 = 4'b1000;
    #200 D3 = 4'b1110;
    #200 D3 = 4'b1000;
    #200 D3 = 4'b0111;
    #200 D3 = 4'b0001;
    #200 D3 = 4'b1110;
    #200 D3 = 4'b1001;
    #200 D3 = 4'b0100;
    #200 D3 = 4'b1111;
    #200 D3 = 4'b0100;
    #200 D3 = 4'b1101;
    #200 D3 = 4'b1111;
    #200 D3 = 4'b0100;
    #200 D3 = 4'b1011;
    #200 D3 = 4'b1100;
    #200 D3 = 4'b1101;
    #200 D3 = 4'b1100;
    #200 D3 = 4'b0110;
    #200 D3 = 4'b1111;
    #200 D3 = 4'b0011;
    #200 D3 = 4'b0001;
    #200 D3 = 4'b1100;
  end

  initial
  begin
    S0 = 1'b0;
    #100 S0 = 1'b1;
    #500 S0 = 1'b0;
    #1400 S0 = 1'b1;
    #900 S0 = 1'b0;
  end

  initial
  begin
    S1 = 1'b0;
    #1000 S1 = 1'b1;
    #600 S1 = 1'b0;
    #600 S1 = 1'b1;
    #400 S1 = 1'b0;
  end

endmodule
