module Accumulator_tb;

reg CLK;
reg Ce;
reg [11:0] Din;
wire [11:0] Dout;
reg RST;

Accumulator
 U0 (
  .CLK(CLK),
  .Ce(Ce),
  .Din(Din),
  .Dout(Dout),
  .RST(RST));

  initial
  begin
    CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
  end

  initial
  begin
    Ce = 1'b1;
  end

  initial
  begin
    Din = 12'b010010000000;
    #200 Din = 12'b100101011100;
    #200 Din = 12'b000100010110;
    #200 Din = 12'b110001010111;
    #200 Din = 12'b110111110100;
    #200 Din = 12'b101111100111;
    #200 Din = 12'b100111110010;
    #200 Din = 12'b100110000100;
    #200 Din = 12'b011100001101;
    #200 Din = 12'b010011000001;
    #200 Din = 12'b010010011100;
    #200 Din = 12'b011110111100;
    #200 Din = 12'b000110111101;
    #200 Din = 12'b101001001000;
    #200 Din = 12'b111010011001;
    #200 Din = 12'b000011010010;
    #200 Din = 12'b011011100001;
    #200 Din = 12'b111101001101;
    #200 Din = 12'b000000000101;
    #200 Din = 12'b110011101110;
    #200 Din = 12'b011001111010;
    #200 Din = 12'b010100010111;
    #200 Din = 12'b001000100010;
    #200 Din = 12'b010000101111;
    #200 Din = 12'b001100000001;
    #200 Din = 12'b110100001011;
    #200 Din = 12'b001000011001;
    #200 Din = 12'b100111111111;
    #200 Din = 12'b111000010110;
    #200 Din = 12'b110100110111;
    #200 Din = 12'b010101111100;
    #200 Din = 12'b100011011001;
    #200 Din = 12'b011100011001;
    #200 Din = 12'b111100110011;
    #200 Din = 12'b000110110001;
    #200 Din = 12'b110010000011;
    #200 Din = 12'b000110010001;
    #200 Din = 12'b100001011101;
    #200 Din = 12'b100011010010;
    #200 Din = 12'b111010100011;
    #200 Din = 12'b000001110010;
    #200 Din = 12'b000110101110;
    #200 Din = 12'b111011001111;
    #200 Din = 12'b010000111110;
    #200 Din = 12'b000100011100;
    #200 Din = 12'b011100111111;
    #200 Din = 12'b001010100010;
    #200 Din = 12'b111010100001;
    #200 Din = 12'b000010101001;
    #200 Din = 12'b010101101010;
  end

  initial
  begin
    RST = 1'b1;
    #200 RST = 1'b0;
  end

endmodule
