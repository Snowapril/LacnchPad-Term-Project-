module MUX4bit_16_tb;

wire [3:0] Dout;
reg S0;
reg S1;
reg S2;
reg S3;
reg [3:0] p0;
reg [3:0] p1;
reg [3:0] p10;
reg [3:0] p11;
reg [3:0] p12;
reg [3:0] p13;
reg [3:0] p14;
reg [3:0] p15;
reg [3:0] p2;
reg [3:0] p3;
reg [3:0] p4;
reg [3:0] p5;
reg [3:0] p6;
reg [3:0] p7;
reg [3:0] p8;
reg [3:0] p9;

MUX4bit_16
 U0 (
  .Dout(Dout),
  .S0(S0),
  .S1(S1),
  .S2(S2),
  .S3(S3),
  .p0(p0),
  .p1(p1),
  .p10(p10),
  .p11(p11),
  .p12(p12),
  .p13(p13),
  .p14(p14),
  .p15(p15),
  .p2(p2),
  .p3(p3),
  .p4(p4),
  .p5(p5),
  .p6(p6),
  .p7(p7),
  .p8(p8),
  .p9(p9));

  initial
  begin
    S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
    #200 S0 = 1'b0;
    #200 S0 = 1'b1;
  end

  initial
  begin
    S1 = 1'b0;
    #400 S1 = 1'b1;
    #400 S1 = 1'b0;
    #400 S1 = 1'b1;
    #400 S1 = 1'b0;
    #400 S1 = 1'b1;
    #400 S1 = 1'b0;
    #400 S1 = 1'b1;
    #400 S1 = 1'b0;
  end

  initial
  begin
    S2 = 1'b0;
    #800 S2 = 1'b1;
    #800 S2 = 1'b0;
    #800 S2 = 1'b1;
  end

  initial
  begin
    S3 = 1'b0;
    #1600 S3 = 1'b1;
  end

  initial
  begin
    p0 = 4'b0101;
    #400 p0 = 4'b0111;
    #200 p0 = 4'b0001;
    #200 p0 = 4'b0101;
    #200 p0 = 4'b1101;
    #200 p0 = 4'b0011;
    #200 p0 = 4'b0010;
    #200 p0 = 4'b0100;
    #200 p0 = 4'b0001;
    #200 p0 = 4'b1001;
    #200 p0 = 4'b1011;
    #200 p0 = 4'b0010;
    #200 p0 = 4'b1101;
    #200 p0 = 4'b0011;
    #200 p0 = 4'b1011;
    #200 p0 = 4'b1101;
    #200 p0 = 4'b0111;
    #200 p0 = 4'b0001;
    #200 p0 = 4'b0110;
    #200 p0 = 4'b0111;
    #200 p0 = 4'b0010;
    #200 p0 = 4'b1001;
    #200 p0 = 4'b0000;
    #200 p0 = 4'b1100;
    #200 p0 = 4'b0111;
    #200 p0 = 4'b1110;
    #200 p0 = 4'b1001;
    #200 p0 = 4'b1101;
    #200 p0 = 4'b0100;
    #200 p0 = 4'b1110;
    #200 p0 = 4'b0100;
    #200 p0 = 4'b1111;
    #200 p0 = 4'b0000;
    #200 p0 = 4'b1110;
    #200 p0 = 4'b1000;
    #200 p0 = 4'b1001;
    #200 p0 = 4'b1110;
    #200 p0 = 4'b0101;
    #200 p0 = 4'b0000;
    #200 p0 = 4'b1000;
    #200 p0 = 4'b0110;
    #200 p0 = 4'b1011;
    #200 p0 = 4'b1101;
    #200 p0 = 4'b0101;
    #200 p0 = 4'b0011;
    #200 p0 = 4'b1100;
    #200 p0 = 4'b0010;
    #400 p0 = 4'b0110;
  end

  initial
  begin
    p1 = 4'b1010;
    #200 p1 = 4'b1011;
    #200 p1 = 4'b0101;
    #200 p1 = 4'b1101;
    #200 p1 = 4'b0011;
    #200 p1 = 4'b1100;
    #200 p1 = 4'b0100;
    #200 p1 = 4'b1110;
    #200 p1 = 4'b0101;
    #200 p1 = 4'b1100;
    #200 p1 = 4'b0101;
    #200 p1 = 4'b0001;
    #200 p1 = 4'b0111;
    #200 p1 = 4'b0110;
    #200 p1 = 4'b1001;
    #200 p1 = 4'b1000;
    #200 p1 = 4'b0111;
    #200 p1 = 4'b1011;
    #200 p1 = 4'b0110;
    #200 p1 = 4'b0101;
    #200 p1 = 4'b0001;
    #200 p1 = 4'b0000;
    #200 p1 = 4'b0101;
    #200 p1 = 4'b1011;
    #200 p1 = 4'b1001;
    #200 p1 = 4'b0000;
    #200 p1 = 4'b1000;
    #200 p1 = 4'b0000;
    #200 p1 = 4'b0010;
    #200 p1 = 4'b1010;
    #200 p1 = 4'b0011;
    #200 p1 = 4'b0101;
    #200 p1 = 4'b1110;
    #200 p1 = 4'b0110;
    #200 p1 = 4'b0001;
    #200 p1 = 4'b0110;
    #200 p1 = 4'b1111;
    #200 p1 = 4'b1001;
    #200 p1 = 4'b1011;
    #200 p1 = 4'b0010;
    #200 p1 = 4'b1011;
    #400 p1 = 4'b1001;
    #200 p1 = 4'b1010;
    #200 p1 = 4'b1111;
    #200 p1 = 4'b0110;
    #200 p1 = 4'b1001;
    #200 p1 = 4'b1110;
    #200 p1 = 4'b0011;
    #200 p1 = 4'b1101;
  end

  initial
  begin
    p10 = 4'b1111;
    #200 p10 = 4'b0000;
    #200 p10 = 4'b0101;
    #200 p10 = 4'b0010;
    #200 p10 = 4'b1111;
    #200 p10 = 4'b0111;
    #200 p10 = 4'b1001;
    #200 p10 = 4'b1101;
    #200 p10 = 4'b0110;
    #200 p10 = 4'b0011;
    #200 p10 = 4'b0101;
    #200 p10 = 4'b1111;
    #200 p10 = 4'b1001;
    #200 p10 = 4'b1011;
    #200 p10 = 4'b1101;
    #400 p10 = 4'b0001;
    #200 p10 = 4'b0011;
    #200 p10 = 4'b1010;
    #200 p10 = 4'b1101;
    #200 p10 = 4'b1011;
    #200 p10 = 4'b1111;
    #200 p10 = 4'b1100;
    #400 p10 = 4'b1101;
    #200 p10 = 4'b0001;
    #200 p10 = 4'b0011;
    #200 p10 = 4'b0000;
    #400 p10 = 4'b1010;
    #200 p10 = 4'b1111;
    #200 p10 = 4'b0111;
    #200 p10 = 4'b0010;
    #200 p10 = 4'b0100;
    #200 p10 = 4'b0000;
    #200 p10 = 4'b0100;
    #200 p10 = 4'b1000;
    #200 p10 = 4'b0100;
    #200 p10 = 4'b0011;
    #200 p10 = 4'b1001;
    #200 p10 = 4'b1000;
    #200 p10 = 4'b1100;
    #200 p10 = 4'b1001;
    #200 p10 = 4'b0011;
    #200 p10 = 4'b0001;
    #200 p10 = 4'b0000;
    #200 p10 = 4'b1001;
    #200 p10 = 4'b0111;
    #200 p10 = 4'b0100;
    #200 p10 = 4'b0001;
  end

  initial
  begin
    p11 = 4'b0001;
    #200 p11 = 4'b0101;
    #200 p11 = 4'b1101;
    #200 p11 = 4'b1010;
    #200 p11 = 4'b1100;
    #200 p11 = 4'b0010;
    #200 p11 = 4'b1111;
    #200 p11 = 4'b1001;
    #200 p11 = 4'b1100;
    #200 p11 = 4'b0001;
    #200 p11 = 4'b1101;
    #200 p11 = 4'b1100;
    #200 p11 = 4'b1101;
    #400 p11 = 4'b1011;
    #200 p11 = 4'b0001;
    #200 p11 = 4'b0111;
    #200 p11 = 4'b1001;
    #200 p11 = 4'b0100;
    #200 p11 = 4'b0111;
    #200 p11 = 4'b0011;
    #200 p11 = 4'b1000;
    #200 p11 = 4'b1111;
    #200 p11 = 4'b1100;
    #200 p11 = 4'b1101;
    #200 p11 = 4'b0000;
    #200 p11 = 4'b0111;
    #200 p11 = 4'b0101;
    #200 p11 = 4'b0000;
    #200 p11 = 4'b0010;
    #200 p11 = 4'b0100;
    #200 p11 = 4'b0001;
    #200 p11 = 4'b0101;
    #400 p11 = 4'b0011;
    #200 p11 = 4'b1111;
    #400 p11 = 4'b1001;
    #200 p11 = 4'b1000;
    #200 p11 = 4'b0101;
    #200 p11 = 4'b0001;
    #400 p11 = 4'b0010;
    #200 p11 = 4'b0011;
    #200 p11 = 4'b0100;
    #200 p11 = 4'b0110;
    #200 p11 = 4'b1001;
    #200 p11 = 4'b0111;
    #200 p11 = 4'b1001;
    #200 p11 = 4'b0101;
  end

  initial
  begin
    p12 = 4'b0011;
    #200 p12 = 4'b1110;
    #200 p12 = 4'b0001;
    #200 p12 = 4'b1000;
    #200 p12 = 4'b1110;
    #200 p12 = 4'b1010;
    #400 p12 = 4'b0011;
    #200 p12 = 4'b0110;
    #400 p12 = 4'b0010;
    #200 p12 = 4'b0111;
    #200 p12 = 4'b0011;
    #200 p12 = 4'b1101;
    #200 p12 = 4'b0000;
    #200 p12 = 4'b0111;
    #200 p12 = 4'b0001;
    #200 p12 = 4'b1011;
    #200 p12 = 4'b0000;
    #200 p12 = 4'b1101;
    #200 p12 = 4'b1110;
    #200 p12 = 4'b0100;
    #200 p12 = 4'b1101;
    #200 p12 = 4'b1100;
    #200 p12 = 4'b0111;
    #200 p12 = 4'b1110;
    #200 p12 = 4'b1011;
    #200 p12 = 4'b1100;
    #400 p12 = 4'b0100;
    #200 p12 = 4'b0101;
    #200 p12 = 4'b0111;
    #200 p12 = 4'b1111;
    #200 p12 = 4'b0011;
    #200 p12 = 4'b1000;
    #200 p12 = 4'b0001;
    #200 p12 = 4'b1011;
    #200 p12 = 4'b0111;
    #200 p12 = 4'b0001;
    #200 p12 = 4'b1011;
    #200 p12 = 4'b0100;
    #400 p12 = 4'b0011;
    #200 p12 = 4'b1111;
    #200 p12 = 4'b1110;
    #200 p12 = 4'b1100;
    #200 p12 = 4'b0001;
    #400 p12 = 4'b1011;
    #200 p12 = 4'b0010;
  end

  initial
  begin
    p13 = 4'b1011;
    #200 p13 = 4'b1001;
    #200 p13 = 4'b1100;
    #200 p13 = 4'b0110;
    #200 p13 = 4'b0101;
    #200 p13 = 4'b1011;
    #200 p13 = 4'b0100;
    #400 p13 = 4'b0111;
    #200 p13 = 4'b0000;
    #200 p13 = 4'b0010;
    #200 p13 = 4'b0011;
    #200 p13 = 4'b1000;
    #200 p13 = 4'b0110;
    #200 p13 = 4'b1010;
    #600 p13 = 4'b0101;
    #400 p13 = 4'b0011;
    #200 p13 = 4'b1111;
    #200 p13 = 4'b0111;
    #400 p13 = 4'b0001;
    #200 p13 = 4'b1011;
    #200 p13 = 4'b1010;
    #200 p13 = 4'b0000;
    #200 p13 = 4'b0100;
    #200 p13 = 4'b1110;
    #200 p13 = 4'b1101;
    #200 p13 = 4'b0000;
    #200 p13 = 4'b1100;
    #200 p13 = 4'b0001;
    #200 p13 = 4'b0000;
    #200 p13 = 4'b1101;
    #200 p13 = 4'b1010;
    #200 p13 = 4'b0001;
    #200 p13 = 4'b1011;
    #200 p13 = 4'b1111;
    #200 p13 = 4'b0000;
    #200 p13 = 4'b0011;
    #200 p13 = 4'b0010;
    #600 p13 = 4'b1010;
    #200 p13 = 4'b0011;
    #200 p13 = 4'b1100;
    #200 p13 = 4'b0100;
    #200 p13 = 4'b0101;
    #200 p13 = 4'b1001;
  end

  initial
  begin
    p14 = 4'b0001;
    #200 p14 = 4'b0111;
    #200 p14 = 4'b1110;
    #200 p14 = 4'b0001;
    #200 p14 = 4'b0011;
    #200 p14 = 4'b1110;
    #200 p14 = 4'b1001;
    #200 p14 = 4'b1000;
    #200 p14 = 4'b0110;
    #200 p14 = 4'b0101;
    #200 p14 = 4'b0100;
    #200 p14 = 4'b1110;
    #200 p14 = 4'b1100;
    #200 p14 = 4'b1010;
    #200 p14 = 4'b0101;
    #200 p14 = 4'b0001;
    #200 p14 = 4'b0101;
    #200 p14 = 4'b1001;
    #200 p14 = 4'b1010;
    #200 p14 = 4'b1110;
    #200 p14 = 4'b1011;
    #200 p14 = 4'b1101;
    #200 p14 = 4'b0100;
    #200 p14 = 4'b0110;
    #200 p14 = 4'b0111;
    #200 p14 = 4'b1011;
    #200 p14 = 4'b0111;
    #200 p14 = 4'b1111;
    #200 p14 = 4'b1011;
    #200 p14 = 4'b0101;
    #200 p14 = 4'b1011;
    #200 p14 = 4'b1101;
    #200 p14 = 4'b1110;
    #200 p14 = 4'b1010;
    #200 p14 = 4'b0010;
    #200 p14 = 4'b0101;
    #200 p14 = 4'b1110;
    #200 p14 = 4'b1001;
    #200 p14 = 4'b0111;
    #200 p14 = 4'b1011;
    #400 p14 = 4'b1000;
    #200 p14 = 4'b1111;
    #200 p14 = 4'b1101;
    #400 p14 = 4'b0001;
    #200 p14 = 4'b0101;
    #200 p14 = 4'b0001;
    #200 p14 = 4'b0000;
  end

  initial
  begin
    p15 = 4'b1001;
    #200 p15 = 4'b1111;
    #200 p15 = 4'b1001;
    #200 p15 = 4'b1000;
    #200 p15 = 4'b1100;
    #200 p15 = 4'b0010;
    #200 p15 = 4'b1101;
    #200 p15 = 4'b1000;
    #200 p15 = 4'b1101;
    #200 p15 = 4'b0110;
    #200 p15 = 4'b1011;
    #200 p15 = 4'b0011;
    #200 p15 = 4'b0101;
    #200 p15 = 4'b1001;
    #200 p15 = 4'b1111;
    #200 p15 = 4'b1110;
    #200 p15 = 4'b0010;
    #200 p15 = 4'b0101;
    #200 p15 = 4'b1100;
    #200 p15 = 4'b1000;
    #200 p15 = 4'b0000;
    #200 p15 = 4'b0111;
    #200 p15 = 4'b1100;
    #200 p15 = 4'b0011;
    #200 p15 = 4'b0110;
    #200 p15 = 4'b1011;
    #200 p15 = 4'b1101;
    #200 p15 = 4'b0100;
    #200 p15 = 4'b1011;
    #200 p15 = 4'b0000;
    #200 p15 = 4'b0111;
    #400 p15 = 4'b1110;
    #200 p15 = 4'b1111;
    #200 p15 = 4'b1101;
    #200 p15 = 4'b1000;
    #200 p15 = 4'b1101;
    #200 p15 = 4'b1110;
    #200 p15 = 4'b0000;
    #200 p15 = 4'b0010;
    #200 p15 = 4'b1110;
    #200 p15 = 4'b0111;
    #200 p15 = 4'b0001;
    #200 p15 = 4'b0111;
    #200 p15 = 4'b1111;
    #200 p15 = 4'b0001;
    #200 p15 = 4'b1100;
    #200 p15 = 4'b1111;
    #200 p15 = 4'b0101;
    #200 p15 = 4'b1000;
  end

  initial
  begin
    p2 = 4'b0000;
    #200 p2 = 4'b1000;
    #200 p2 = 4'b1101;
    #200 p2 = 4'b0100;
    #400 p2 = 4'b0010;
    #200 p2 = 4'b0011;
    #200 p2 = 4'b1101;
    #200 p2 = 4'b1000;
    #200 p2 = 4'b1101;
    #200 p2 = 4'b0011;
    #400 p2 = 4'b1111;
    #200 p2 = 4'b0101;
    #200 p2 = 4'b1011;
    #200 p2 = 4'b0010;
    #200 p2 = 4'b0100;
    #200 p2 = 4'b1001;
    #200 p2 = 4'b1111;
    #200 p2 = 4'b0101;
    #200 p2 = 4'b1000;
    #200 p2 = 4'b0010;
    #200 p2 = 4'b0001;
    #400 p2 = 4'b1100;
    #400 p2 = 4'b0110;
    #200 p2 = 4'b0111;
    #200 p2 = 4'b1100;
    #200 p2 = 4'b0001;
    #200 p2 = 4'b0100;
    #200 p2 = 4'b1010;
    #200 p2 = 4'b0110;
    #200 p2 = 4'b0000;
    #200 p2 = 4'b0110;
    #200 p2 = 4'b0001;
    #200 p2 = 4'b1010;
    #200 p2 = 4'b0011;
    #200 p2 = 4'b1111;
    #200 p2 = 4'b0011;
    #200 p2 = 4'b0111;
    #200 p2 = 4'b1010;
    #200 p2 = 4'b1111;
    #200 p2 = 4'b1000;
    #200 p2 = 4'b0110;
    #200 p2 = 4'b1010;
    #400 p2 = 4'b0111;
    #200 p2 = 4'b0011;
    #200 p2 = 4'b1001;
  end

  initial
  begin
    p3 = 4'b0001;
    #200 p3 = 4'b1010;
    #200 p3 = 4'b0010;
    #200 p3 = 4'b0110;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b1111;
    #200 p3 = 4'b1100;
    #200 p3 = 4'b0011;
    #200 p3 = 4'b0101;
    #200 p3 = 4'b1110;
    #200 p3 = 4'b0110;
    #200 p3 = 4'b1010;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b1011;
    #200 p3 = 4'b0010;
    #200 p3 = 4'b1011;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b1010;
    #200 p3 = 4'b1111;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b1011;
    #200 p3 = 4'b0111;
    #200 p3 = 4'b1111;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b0010;
    #200 p3 = 4'b0000;
    #200 p3 = 4'b1011;
    #200 p3 = 4'b0000;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b0011;
    #200 p3 = 4'b1110;
    #200 p3 = 4'b0111;
    #200 p3 = 4'b0001;
    #400 p3 = 4'b1111;
    #200 p3 = 4'b0010;
    #400 p3 = 4'b1100;
    #200 p3 = 4'b0111;
    #200 p3 = 4'b1101;
    #400 p3 = 4'b1111;
    #200 p3 = 4'b1010;
    #200 p3 = 4'b1101;
    #200 p3 = 4'b0111;
    #200 p3 = 4'b0011;
    #200 p3 = 4'b0000;
    #200 p3 = 4'b1000;
    #200 p3 = 4'b1010;
    #200 p3 = 4'b0111;
  end

  initial
  begin
    p4 = 4'b1101;
    #200 p4 = 4'b1010;
    #200 p4 = 4'b1011;
    #200 p4 = 4'b1000;
    #200 p4 = 4'b0100;
    #200 p4 = 4'b0010;
    #200 p4 = 4'b0111;
    #200 p4 = 4'b1000;
    #200 p4 = 4'b0000;
    #200 p4 = 4'b1011;
    #200 p4 = 4'b0011;
    #200 p4 = 4'b1011;
    #200 p4 = 4'b1110;
    #200 p4 = 4'b0110;
    #200 p4 = 4'b0011;
    #200 p4 = 4'b0110;
    #200 p4 = 4'b1101;
    #200 p4 = 4'b1011;
    #200 p4 = 4'b0000;
    #200 p4 = 4'b1011;
    #200 p4 = 4'b0001;
    #200 p4 = 4'b1100;
    #200 p4 = 4'b1001;
    #200 p4 = 4'b1010;
    #200 p4 = 4'b1101;
    #200 p4 = 4'b0110;
    #200 p4 = 4'b0111;
    #200 p4 = 4'b1011;
    #200 p4 = 4'b1100;
    #200 p4 = 4'b0000;
    #200 p4 = 4'b0111;
    #400 p4 = 4'b0011;
    #200 p4 = 4'b1010;
    #200 p4 = 4'b0100;
    #200 p4 = 4'b0000;
    #200 p4 = 4'b1110;
    #200 p4 = 4'b0111;
    #200 p4 = 4'b0101;
    #200 p4 = 4'b0011;
    #200 p4 = 4'b1111;
    #200 p4 = 4'b0010;
    #200 p4 = 4'b1001;
    #200 p4 = 4'b0100;
    #200 p4 = 4'b0111;
    #200 p4 = 4'b0100;
    #200 p4 = 4'b1001;
    #200 p4 = 4'b1110;
    #200 p4 = 4'b0000;
    #200 p4 = 4'b0101;
  end

  initial
  begin
    p5 = 4'b0100;
    #200 p5 = 4'b1010;
    #200 p5 = 4'b0111;
    #200 p5 = 4'b0000;
    #200 p5 = 4'b0111;
    #400 p5 = 4'b0101;
    #200 p5 = 4'b1011;
    #200 p5 = 4'b0000;
    #400 p5 = 4'b0100;
    #400 p5 = 4'b0011;
    #200 p5 = 4'b1110;
    #200 p5 = 4'b0111;
    #200 p5 = 4'b0010;
    #200 p5 = 4'b0011;
    #200 p5 = 4'b1111;
    #200 p5 = 4'b1001;
    #200 p5 = 4'b1010;
    #200 p5 = 4'b0010;
    #200 p5 = 4'b1100;
    #200 p5 = 4'b0000;
    #200 p5 = 4'b1110;
    #200 p5 = 4'b0000;
    #200 p5 = 4'b0110;
    #200 p5 = 4'b1111;
    #200 p5 = 4'b0100;
    #200 p5 = 4'b0110;
    #200 p5 = 4'b0111;
    #200 p5 = 4'b1001;
    #200 p5 = 4'b0001;
    #400 p5 = 4'b0011;
    #200 p5 = 4'b0101;
    #200 p5 = 4'b0100;
    #200 p5 = 4'b0110;
    #200 p5 = 4'b1011;
    #200 p5 = 4'b1110;
    #200 p5 = 4'b0010;
    #200 p5 = 4'b1100;
    #200 p5 = 4'b0000;
    #200 p5 = 4'b1110;
    #200 p5 = 4'b1011;
    #200 p5 = 4'b0001;
    #200 p5 = 4'b0110;
    #200 p5 = 4'b0101;
    #200 p5 = 4'b1010;
    #200 p5 = 4'b0110;
    #200 p5 = 4'b1110;
  end

  initial
  begin
    p6 = 4'b0100;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b1010;
    #200 p6 = 4'b0010;
    #200 p6 = 4'b1010;
    #200 p6 = 4'b0001;
    #200 p6 = 4'b0010;
    #200 p6 = 4'b0011;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b1110;
    #200 p6 = 4'b0010;
    #200 p6 = 4'b1010;
    #200 p6 = 4'b1000;
    #200 p6 = 4'b0011;
    #200 p6 = 4'b1001;
    #200 p6 = 4'b0010;
    #200 p6 = 4'b1000;
    #200 p6 = 4'b0101;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b0001;
    #200 p6 = 4'b1000;
    #200 p6 = 4'b1010;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b0010;
    #200 p6 = 4'b0110;
    #200 p6 = 4'b1100;
    #200 p6 = 4'b1010;
    #200 p6 = 4'b0111;
    #200 p6 = 4'b0001;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b0011;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b0110;
    #200 p6 = 4'b0101;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b0111;
    #200 p6 = 4'b1101;
    #200 p6 = 4'b0100;
    #600 p6 = 4'b0001;
    #200 p6 = 4'b0110;
    #200 p6 = 4'b0101;
    #200 p6 = 4'b0011;
    #200 p6 = 4'b1001;
    #200 p6 = 4'b0001;
    #200 p6 = 4'b0010;
    #200 p6 = 4'b0111;
    #400 p6 = 4'b0101;
  end

  initial
  begin
    p7 = 4'b1111;
    #200 p7 = 4'b1110;
    #200 p7 = 4'b1010;
    #200 p7 = 4'b1001;
    #200 p7 = 4'b0000;
    #200 p7 = 4'b0001;
    #200 p7 = 4'b1010;
    #200 p7 = 4'b0010;
    #200 p7 = 4'b0011;
    #200 p7 = 4'b0010;
    #200 p7 = 4'b1111;
    #200 p7 = 4'b0001;
    #200 p7 = 4'b1100;
    #200 p7 = 4'b0011;
    #200 p7 = 4'b1111;
    #200 p7 = 4'b0001;
    #200 p7 = 4'b1010;
    #200 p7 = 4'b0000;
    #200 p7 = 4'b1110;
    #200 p7 = 4'b1011;
    #200 p7 = 4'b1010;
    #400 p7 = 4'b0010;
    #200 p7 = 4'b0000;
    #200 p7 = 4'b0011;
    #200 p7 = 4'b1011;
    #200 p7 = 4'b0110;
    #200 p7 = 4'b1001;
    #200 p7 = 4'b0101;
    #200 p7 = 4'b0000;
    #200 p7 = 4'b0110;
    #200 p7 = 4'b1101;
    #200 p7 = 4'b1111;
    #400 p7 = 4'b1100;
    #200 p7 = 4'b1111;
    #400 p7 = 4'b1110;
    #200 p7 = 4'b0001;
    #200 p7 = 4'b0101;
    #400 p7 = 4'b1010;
    #200 p7 = 4'b0100;
    #200 p7 = 4'b1010;
    #200 p7 = 4'b0110;
    #200 p7 = 4'b0010;
    #200 p7 = 4'b0101;
    #200 p7 = 4'b1100;
    #200 p7 = 4'b0011;
    #200 p7 = 4'b0001;
  end

  initial
  begin
    p8 = 4'b0011;
    #400 p8 = 4'b0111;
    #200 p8 = 4'b0010;
    #200 p8 = 4'b1010;
    #200 p8 = 4'b1100;
    #200 p8 = 4'b1000;
    #200 p8 = 4'b0001;
    #200 p8 = 4'b0111;
    #200 p8 = 4'b0011;
    #200 p8 = 4'b0110;
    #200 p8 = 4'b0111;
    #200 p8 = 4'b1110;
    #200 p8 = 4'b0000;
    #200 p8 = 4'b0101;
    #600 p8 = 4'b1000;
    #200 p8 = 4'b0101;
    #200 p8 = 4'b0011;
    #200 p8 = 4'b0110;
    #200 p8 = 4'b1101;
    #200 p8 = 4'b1100;
    #200 p8 = 4'b1010;
    #200 p8 = 4'b0001;
    #400 p8 = 4'b1101;
    #200 p8 = 4'b1110;
    #400 p8 = 4'b0110;
    #200 p8 = 4'b0111;
    #200 p8 = 4'b0001;
    #200 p8 = 4'b1000;
    #200 p8 = 4'b0011;
    #200 p8 = 4'b0001;
    #400 p8 = 4'b1111;
    #200 p8 = 4'b0001;
    #200 p8 = 4'b0011;
    #200 p8 = 4'b0111;
    #200 p8 = 4'b1101;
    #200 p8 = 4'b0000;
    #200 p8 = 4'b0011;
    #200 p8 = 4'b0111;
    #200 p8 = 4'b1110;
    #200 p8 = 4'b1010;
    #200 p8 = 4'b0010;
    #200 p8 = 4'b0101;
    #200 p8 = 4'b1111;
    #200 p8 = 4'b0101;
  end

  initial
  begin
    p9 = 4'b0110;
    #200 p9 = 4'b0010;
    #200 p9 = 4'b0011;
    #200 p9 = 4'b0100;
    #200 p9 = 4'b1010;
    #200 p9 = 4'b1011;
    #200 p9 = 4'b1111;
    #200 p9 = 4'b1001;
    #200 p9 = 4'b1111;
    #200 p9 = 4'b0011;
    #200 p9 = 4'b0001;
    #200 p9 = 4'b0100;
    #200 p9 = 4'b0001;
    #200 p9 = 4'b0000;
    #200 p9 = 4'b1111;
    #200 p9 = 4'b0010;
    #200 p9 = 4'b0000;
    #200 p9 = 4'b0110;
    #200 p9 = 4'b1000;
    #400 p9 = 4'b0000;
    #200 p9 = 4'b0010;
    #200 p9 = 4'b0000;
    #200 p9 = 4'b0100;
    #200 p9 = 4'b1001;
    #200 p9 = 4'b0101;
    #200 p9 = 4'b0000;
    #200 p9 = 4'b0101;
    #200 p9 = 4'b1111;
    #200 p9 = 4'b0100;
    #200 p9 = 4'b1000;
    #200 p9 = 4'b0000;
    #200 p9 = 4'b0100;
    #200 p9 = 4'b1010;
    #200 p9 = 4'b0001;
    #200 p9 = 4'b0100;
    #200 p9 = 4'b0010;
    #200 p9 = 4'b1110;
    #200 p9 = 4'b1011;
    #200 p9 = 4'b0111;
    #200 p9 = 4'b1110;
    #200 p9 = 4'b0111;
    #200 p9 = 4'b1010;
    #200 p9 = 4'b0010;
    #400 p9 = 4'b0000;
    #200 p9 = 4'b1111;
    #200 p9 = 4'b1110;
    #200 p9 = 4'b1011;
    #200 p9 = 4'b0101;
  end

endmodule
